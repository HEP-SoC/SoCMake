module top;

 mod1 mod1_i();

endmodule;
