`define INCLUDED_NUM 55
