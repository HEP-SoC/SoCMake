module mod1;

    submod1 submod1_i();

endmodule;
