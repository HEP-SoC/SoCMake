module tb;
 initial begin
     $display("Simulated with Iverilog, from SoCMake build system\n");
     $finish();
 end
 endmodule
