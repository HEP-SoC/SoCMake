module submod1;

endmodule;

