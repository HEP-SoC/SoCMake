module top1;
    initial begin
        $display("Module top1\n");
        $fatal();
    end
endmodule
