module top2;
    initial begin
        $display("Module top2\n");
        $finish();
    end
endmodule

