module submod2;

endmodule;


