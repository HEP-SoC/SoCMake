module tb;
 initial begin
     $display("Hello world, from SoCMake build system\n");
     $finish();
 end
 endmodule
