module tb;

 printer_0 printer_0_i ();
 printer_1 printer_1_i ();
 printer_2 printer_2_i ();
 printer_3 printer_3_i ();
 printer_4 printer_4_i ();
 printer_5 printer_5_i ();
 printer_6 printer_6_i ();
 printer_7 printer_7_i ();
 printer_8 printer_8_i ();
 printer_9 printer_9_i ();
 printer_10 printer_10_i ();
 printer_11 printer_11_i ();
 printer_12 printer_12_i ();
 printer_13 printer_13_i ();
 printer_14 printer_14_i ();
 printer_15 printer_15_i ();
 printer_16 printer_16_i ();
 printer_17 printer_17_i ();
 printer_18 printer_18_i ();
 printer_19 printer_19_i ();
 printer_20 printer_20_i ();
 printer_21 printer_21_i ();
 printer_22 printer_22_i ();
 printer_23 printer_23_i ();
 printer_24 printer_24_i ();
 printer_25 printer_25_i ();
 printer_26 printer_26_i ();
 printer_27 printer_27_i ();
 printer_28 printer_28_i ();
 printer_29 printer_29_i ();
 printer_30 printer_30_i ();
 printer_31 printer_31_i ();
 printer_32 printer_32_i ();

 initial begin
     $display("Hello world, from SoCMake build system\n");
     $finish();
 end
 endmodule
